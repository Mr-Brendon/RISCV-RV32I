--Il PC per le istruzioni normali si incrementa di 4 perche sono lunghe 4 byte ciascuna (quelle normali).

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity PC is
    port(CLK: in std_logic;
         
         );
end PC;

architecture PC_bh of PC is

begin


end PC_bh;
