----------------------------------------------------------------------------------
-- Engineer: 
-- 
-- Create Date: 13.11.2024
-- Module Name: RISCV_Core
-- Project Name: RISCV CPU RV32I instruction set
--
-- Description:
--

----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;
--library UNISIM;
--use UNISIM.VComponents.all;

entity RISCV_Core is
end RISCV_Core;

architecture Core of RISCV_Core is

begin


end Core;
