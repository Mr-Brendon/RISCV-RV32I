
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package Instruments_pkg is
--Constants:
constant Nbit: integer := 32;
constant binary4in32: std_logic_vector(31 downto 0) := "00000000000000000000000000000100";
end Instruments_pkg;
